module or_dut (
    input a,b ,output y
);

or(y,a,b);
// assign y=a^b;
    
endmodule
 