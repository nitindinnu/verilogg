module serial_adder (
    
);

endmodule //serial_adder
