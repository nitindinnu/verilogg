module and_tb_param (
);
    reg [n-1:0]a,b;
    output y;  

    and_dut_param a1(y,a,b);
    initial begin
        
    end
endmodule
