module  ha(input a,b,output y,c);
assign y= a^b;
assign c=a&b;   
endmodule
