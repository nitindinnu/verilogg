module xor_dut (
    input a,b,c,d ,output y
);

xor(y,a,b,c,d);
// assign y=a^b;
    
endmodule
 
