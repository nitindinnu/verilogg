module dec_to_bin (
    input dec,output bin
);
    integer dec = 3'd8;
    $display("binary is =%0d",dec);
endmodule
