module mux8x1_using_4x1_dut (
    i,s,y
);
  input [0:7]i;  
  input [2:0]s;  
  output [2:0]y;

  assign y[0]=s[0]? (s[1]?i[3]:i[2]) : (s[1]?i[1]:i[0]);
  assign y[1]=s[0]? (s[1]?i[7]:i[6]) : (s[1]?i[5]:i[4]);
  
  assign y[2]=s[2]?y[1]:y[0];

endmodule

module mux8x1_using_4x1_tb (
    
);
    reg [0:7]i;  
    reg [2:0]s;  
    wire [2:0]y;

mux8x1_using_4x1_dut ab(i,s,y);
    initial begin
        #10;
        s[2]=0;s[1]=0;s[0]=0;  i[0]=1;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=0; #10;
        s[2]=0;s[1]=0;s[0]=1;  i[0]=0;i[1]=1;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=0; #10;
        s[2]=0;s[1]=1;s[0]=0;  i[0]=0;i[1]=0;i[2]=1;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=0; #10;
        s[2]=0;s[1]=1;s[0]=1;  i[0]=0;i[1]=0;i[2]=0;i[3]=1;i[4]=0;i[5]=0;i[6]=0;i[7]=0; #10;
        s[2]=1;s[1]=0;s[0]=0;  i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=1;i[5]=0;i[6]=0;i[7]=0; #10;
        s[2]=1;s[1]=0;s[0]=1;  i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=1;i[6]=0;i[7]=0; #10;
        s[2]=1;s[1]=1;s[0]=0;  i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=1;i[7]=0; #10;
        s[2]=1;s[1]=1;s[0]=1;  i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=1; #10;
    end
endmodule

